module REDUCTION1(
  input [25:0]pp0, pp1, pp2, pp3, pp4, pp5, pp6, pp7, pp8, pp9, pp10,
  input [24:0]pp11,
  input [22:0]pp12,
  
  output [47:0]red1_0,
  output [44:0]red1_1,
  output [41:0]red1_2,
  output [37:0]red1_3,
  output [33:0]red1_4,
  output [29:0]red1_5,
  output [25:0]red1_6,
  output [21:0]red1_7,
  output [17:0]red1_8,
  output [13:0]red1_9,
  output [9:0]red1_10,
  output [5:0]red1_11,
  output [1:0]red1_12);
  
  half half1_0[9:0](
    .A({pp0[21], pp0[19], pp0[17], pp0[15], pp0[13], pp0[11], pp0[9], pp0[7], pp0[5], pp0[3]}),
    .B({pp1[19], pp1[17], pp1[15], pp1[13], pp1[11], pp1[9], pp1[7], pp1[5], pp1[3], pp1[1]}),
    .S({red1_0[21], red1_0[19], red1_0[17], red1_0[15], red1_0[13], red1_0[11], red1_0[9], red1_0[7], red1_0[5], red1_0[3]}),
    .Cout({red1_0[22], red1_0[20], red1_0[18], red1_0[16], red1_0[14], red1_0[12], red1_0[10], red1_0[8], red1_0[6], red1_0[4]}));
  
  assign red1_0[23] = !pp0[23];
  assign red1_0[24] = pp0[23];
  
  assign red1_0[47:25] = {
    pp11[24:23],
    pp10[25:24],
    pp9[25:24],
    pp8[25:24],
    pp7[25:24],
    pp6[25:24],
    pp5[25:24],
    pp4[25:24],
    pp3[25:24],
    pp2[25:24],
    pp1[25:24],
    pp0[25]};
  assign red1_0[2:0] = pp0[2:0];
  
  assign red1_1[44:0] = {
    pp12[22:21],
    pp11[22:21],
    pp10[23:22],
    pp9[23:22],
    pp8[23:22],
    pp7[23:22],
    pp6[23:22],
    pp5[23:22],
    pp4[23:22],
    pp3[23:22],
    pp2[23:22],
    pp1[23],
    pp0[24], pp1[21],
    pp0[22], pp2[17],
    pp0[20], pp2[15],
    pp0[18], pp2[13],
    pp0[16], pp2[11],
    pp0[14], pp2[9],
    pp0[12], pp2[7],
    pp0[10],  pp2[5],
    pp0[8],  pp2[3],
    pp0[6],  pp2[1],
    pp0[4],  pp1[0]};
  
  assign red1_2[41:0] = {
    pp12[20:19],
    pp11[20:19],
    pp10[21:20],
    pp9[21:20],
    pp8[21:20],
    pp7[21:20],
    pp6[21:20],
    pp5[21:20],
    pp4[21:20],
    pp3[21:20],
    pp2[21],
    pp1[22], pp2[19],
    pp1[20], pp3[15],
    pp1[18], pp3[13],
    pp1[16], pp3[11],
    pp1[14], pp3[9],
    pp1[12], pp3[7],
    pp1[10], pp3[5],
    pp1[8],  pp3[3],
    pp1[6],  pp3[1],
    pp1[4],  pp2[0],
    pp1[2]};
  
  assign red1_3[37:0] = {
    pp12[18:17],
    pp11[18:17],
    pp10[19:18],
    pp9[19:18],
    pp8[19:18],
    pp7[19:18],
    pp6[19:18],
    pp5[19:18],
    pp4[19:18],
    pp3[19],
    pp2[20], pp3[17],
    pp2[18], pp4[13],
    pp2[16], pp4[11],
    pp2[14], pp4[9],
    pp2[12], pp4[7],
    pp2[10], pp4[5],
    pp2[8],  pp4[3],
    pp2[6],  pp4[1],
    pp2[4],  pp3[0],
    pp2[2]};
  
  assign red1_4[33:0] = {
    pp12[16:15],
    pp11[16:15],
    pp10[17:16],
    pp9[17:16],
    pp8[17:16],
    pp7[17:16],
    pp6[17:16],
    pp5[17:16],
    pp4[17],
    pp3[18], pp4[15],
    pp3[16], pp5[11],
    pp3[14], pp5[9],
    pp3[12], pp5[7],
    pp3[10], pp5[5],
    pp3[8],  pp5[3],
    pp3[6],  pp5[1],
    pp3[4],  pp4[0],
    pp3[2]};
  
  assign red1_5[29:0] = {
    pp12[14:13],
    pp11[14:13],
    pp10[15:14],
    pp9[15:14],
    pp8[15:14],
    pp7[15:14],
    pp6[15:14],
    pp5[15],
    pp4[16], pp5[13],
    pp4[14], pp6[9],
    pp4[12], pp6[7],
    pp4[10], pp6[5],
    pp4[8],  pp6[3],
    pp4[6],  pp6[1],
    pp4[4],  pp5[0],
    pp4[2]};
  
  assign red1_6[25:0] = {
    pp12[12:11],
    pp11[12:11],
    pp10[13:12],
    pp9[13:12],
    pp8[13:12],
    pp7[13:12],
    pp6[13],
    pp5[14], pp6[11],
    pp5[12], pp7[7],
    pp5[10], pp7[5],
    pp5[8],  pp7[3],
    pp5[6],  pp7[1],
    pp5[4],  pp6[0],
    pp5[2]};
  
  assign red1_7[21:0] = {
    pp12[10:9],
    pp11[10:9],
    pp10[11:10],
    pp9[11:10],
    pp8[11:10],
    pp7[11],
    pp6[12], pp7[9],
    pp6[10], pp8[5],
    pp6[8],  pp8[3],
    pp6[6],  pp8[1],
    pp6[4],  pp7[0],
    pp6[2]};
  
  assign red1_8[17:0] = {
    pp12[8:7],
    pp11[8:7],
    pp10[9:8],
    pp9[9:8],
    pp8[9],
    pp7[10], pp8[7],
    pp7[8],  pp9[3],
    pp7[6],  pp9[1],
    pp7[4],  pp8[0],
    pp7[2]};
  
  assign red1_9[13:0] = {
    pp12[6:5],
    pp11[6:5],
    pp10[7:6],
    pp9[7],
    pp8[8], pp9[5],
    pp8[6], pp10[1],
    pp8[4], pp9[0],
    pp8[2]};
  
  assign red1_10[9:0] = {
    pp12[4:3],
    pp11[4:3],
    pp10[5],
    pp9[6], pp10[3],
    pp9[4], pp10[0],
    pp9[2]};
  
  assign red1_11[5:0] = {
    pp12[2:1],
    pp11[2],
    pp10[4], pp11[0],
    pp10[2]};
  
  assign red1_12[1:0] = {
    pp12[0],
    pp11[1]};
  
endmodule
