testbench goes here
